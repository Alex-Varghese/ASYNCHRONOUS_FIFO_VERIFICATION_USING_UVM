`define num_of_txns 16

`define DSIZE 8
`define DEPTH 16

`define ASIZE 4

`define test 1 

`define run_all 0 
