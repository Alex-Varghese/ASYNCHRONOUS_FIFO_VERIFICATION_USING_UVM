`define ASIZE 4
`define DSIZE 8
`define no_of_txns 5
