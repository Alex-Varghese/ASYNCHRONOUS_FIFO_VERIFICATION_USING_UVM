
package async_fifo_pkg;

`include "async_fifo_seq_item.sv"
`include "async_fifo_seq_base.sv"
`include "async_fifo_seq_random.sv"

`include "async_fifo_sequencer.sv"
`include "async_fifo_driver.sv"
`include "async_fifo_write_monitor.sv"
`include "async_fifo_read_monitor.sv"
`include "async_fifo_write_agent.sv"
`include "async_fifo_read_agent.sv"
`include "async_fifo_scoreboard.sv"
`include "../coverage/subscriber.sv"
		
endpackage:async_fifo_pkg
