/*
 //coverage start
 covergroup FIFO_coverage;
 	option.per_instance = 1;

  	WRITE_DATA : coverpoint DUV_IF.wdata{
		option.comment = "write data ";
	}


	WDATA_BOUNDARY: coverpoint DUV_IF.wdata {
		option.comment = "boundary write data ";
    		bins wdata_boundary[] = {9'hff,9'h00};

        }


	FULL : coverpoint DUV_IF.wfull {
		option.comment = "FULL_FLAG";
		bins full_c   = { 0  };
		bins full_c1  = { 1  };
	}

	EMPTY: coverpoint DUV_IF.rempty {
		option.comment = "WHEN RESET IS OFF check EMPTY";
		bins empty_c  = {0 };
		bins empty_c1 = {1 };
	}



  	READ_DATA : coverpoint DUV_IF.rdata{
		option.comment = "read data ";
	}

	WRITE_INC : coverpoint DUV_IF.winc{
  		bins incr_s = (0 => 1);
 		bins incr_s1 = (1 => 0);
  	}

  	READ_INC : coverpoint DUV_IF.rinc{
  		bins incr_sr = (0 => 1);
  		bins incr_s1r = (1 => 0);
  	}

	WRITE_CLK: coverpoint DUV_IF.wclk {
  		option.comment = "write clock signal";
  		bins clk_low_to_high = (0 => 1);
  		bins clk_high_to_low = (1 => 0);
	}

	READ_CLK: coverpoint DUV_IF.rclk {
  		option.comment = "read clock signal";
  		bins clk_low_to_high = (0 => 1);
  		bins clk_high_to_low = (1 => 0);
	}

WRITExADDxDATA : cross WRITE_INC,WRITE_DATA;
READxADDxDATA  : cross READ_INC, READ_DATA;
READxWRITE     : cross  WRITE_DATA,READ_DATA;

endgroup


*/
